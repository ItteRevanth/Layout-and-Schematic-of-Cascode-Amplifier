magic
tech scmos
timestamp 1699376808
<< nwell >>
rect -248 -80 -87 82
<< polysilicon >>
rect -109 63 -106 67
rect -110 61 -106 63
rect -110 11 -106 13
rect -110 7 -107 11
rect -231 -13 -228 -9
rect -110 -11 -107 -7
rect -232 -14 -228 -13
rect -191 -14 -187 -11
rect -110 -14 -106 -11
rect -146 -56 -142 -52
rect -232 -64 -228 -62
rect -191 -64 -187 -62
rect -232 -68 -229 -64
rect -190 -68 -187 -64
rect -146 -64 -142 -62
rect -110 -64 -106 -62
rect -146 -68 -143 -64
rect -109 -68 -106 -64
rect -232 -106 -229 -102
rect -190 -106 -187 -102
rect -232 -108 -228 -106
rect -191 -108 -187 -106
rect -146 -106 -143 -102
rect -109 -106 -106 -102
rect -146 -108 -142 -106
rect -110 -108 -106 -106
rect -191 -131 -187 -128
rect -191 -132 -165 -131
rect -146 -131 -142 -128
rect -110 -131 -106 -128
rect -161 -132 -142 -131
rect -191 -135 -142 -132
rect -232 -141 -228 -138
rect -191 -151 -173 -150
rect -169 -151 -143 -150
rect -191 -153 -143 -151
rect -191 -156 -187 -153
rect -146 -154 -143 -153
rect -109 -154 -106 -150
rect -146 -156 -142 -154
rect -110 -156 -106 -154
rect -191 -179 -187 -176
rect -146 -179 -142 -176
rect -110 -179 -106 -176
<< ndiffusion >>
rect -233 -112 -232 -108
rect -237 -138 -232 -112
rect -228 -134 -223 -108
rect -196 -124 -191 -108
rect -192 -128 -191 -124
rect -187 -112 -186 -108
rect -187 -128 -182 -112
rect -147 -112 -146 -108
rect -151 -128 -146 -112
rect -142 -124 -137 -108
rect -142 -128 -141 -124
rect -115 -124 -110 -108
rect -111 -128 -110 -124
rect -106 -112 -105 -108
rect -106 -128 -101 -112
rect -228 -138 -227 -134
rect -192 -160 -191 -156
rect -196 -176 -191 -160
rect -187 -172 -182 -156
rect -187 -176 -186 -172
rect -147 -160 -146 -156
rect -151 -176 -146 -160
rect -142 -172 -137 -156
rect -142 -176 -141 -172
rect -115 -172 -110 -156
rect -111 -176 -110 -172
rect -106 -160 -105 -156
rect -106 -176 -101 -160
<< pdiffusion >>
rect -115 17 -110 61
rect -111 13 -110 17
rect -106 57 -105 61
rect -106 13 -101 57
rect -237 -58 -232 -14
rect -233 -62 -232 -58
rect -228 -18 -227 -14
rect -228 -62 -223 -18
rect -192 -18 -191 -14
rect -196 -62 -191 -18
rect -187 -58 -182 -14
rect -111 -18 -110 -14
rect -187 -62 -186 -58
rect -151 -58 -146 -56
rect -147 -62 -146 -58
rect -142 -60 -141 -56
rect -142 -62 -137 -60
rect -115 -62 -110 -18
rect -106 -58 -101 -14
rect -106 -62 -105 -58
<< metal1 >>
rect -235 72 -227 76
rect -223 72 -196 76
rect -192 72 -166 76
rect -162 72 -141 76
rect -137 72 -123 76
rect -119 72 -105 76
rect -101 72 -94 76
rect -238 -13 -235 -9
rect -227 -14 -223 72
rect -196 -14 -192 72
rect -141 -56 -137 72
rect -119 63 -113 67
rect -105 61 -101 72
rect -115 -14 -111 13
rect -103 7 -92 11
rect -103 -11 -100 -7
rect -237 -87 -233 -62
rect -225 -68 -194 -64
rect -186 -87 -182 -62
rect -151 -83 -147 -62
rect -139 -68 -113 -64
rect -105 -65 -101 -62
rect -96 -65 -92 7
rect -137 -83 -133 -68
rect -151 -87 -133 -83
rect -105 -69 -92 -65
rect -237 -91 -220 -87
rect -237 -108 -233 -91
rect -224 -102 -220 -91
rect -186 -91 -169 -87
rect -225 -106 -194 -102
rect -186 -108 -182 -91
rect -227 -186 -223 -138
rect -196 -156 -192 -128
rect -173 -147 -169 -91
rect -151 -108 -147 -87
rect -139 -106 -113 -102
rect -105 -108 -101 -69
rect -165 -128 -161 -123
rect -141 -139 -137 -128
rect -151 -143 -137 -139
rect -115 -140 -111 -128
rect -151 -156 -147 -143
rect -115 -144 -101 -140
rect -139 -154 -113 -150
rect -105 -156 -101 -144
rect -186 -186 -182 -176
rect -141 -186 -137 -176
rect -115 -186 -111 -176
rect -240 -190 -227 -186
rect -223 -190 -208 -186
rect -204 -190 -186 -186
rect -182 -190 -161 -186
rect -157 -190 -141 -186
rect -137 -190 -115 -186
rect -111 -190 -98 -186
<< ntransistor >>
rect -232 -138 -228 -108
rect -191 -128 -187 -108
rect -146 -128 -142 -108
rect -110 -128 -106 -108
rect -191 -176 -187 -156
rect -146 -176 -142 -156
rect -110 -176 -106 -156
<< ptransistor >>
rect -110 13 -106 61
rect -232 -62 -228 -14
rect -191 -62 -187 -14
rect -146 -62 -142 -56
rect -110 -62 -106 -14
<< polycontact >>
rect -113 63 -109 67
rect -107 7 -103 11
rect -235 -13 -231 -9
rect -107 -11 -103 -7
rect -229 -68 -225 -64
rect -194 -68 -190 -64
rect -143 -68 -139 -64
rect -113 -68 -109 -64
rect -229 -106 -225 -102
rect -194 -106 -190 -102
rect -143 -106 -139 -102
rect -113 -106 -109 -102
rect -165 -132 -161 -128
rect -173 -151 -169 -147
rect -143 -154 -139 -150
rect -113 -154 -109 -150
<< ndcontact >>
rect -237 -112 -233 -108
rect -196 -128 -192 -124
rect -186 -112 -182 -108
rect -151 -112 -147 -108
rect -141 -128 -137 -124
rect -115 -128 -111 -124
rect -105 -112 -101 -108
rect -227 -138 -223 -134
rect -196 -160 -192 -156
rect -186 -176 -182 -172
rect -151 -160 -147 -156
rect -141 -176 -137 -172
rect -115 -176 -111 -172
rect -105 -160 -101 -156
<< pdcontact >>
rect -115 13 -111 17
rect -105 57 -101 61
rect -237 -62 -233 -58
rect -227 -18 -223 -14
rect -196 -18 -192 -14
rect -115 -18 -111 -14
rect -186 -62 -182 -58
rect -151 -62 -147 -58
rect -141 -60 -137 -56
rect -105 -62 -101 -58
<< psubstratepcontact >>
rect -244 -190 -240 -186
rect -227 -190 -223 -186
rect -208 -190 -204 -186
rect -186 -190 -182 -186
rect -161 -190 -157 -186
rect -141 -190 -137 -186
rect -115 -190 -111 -186
rect -98 -190 -94 -186
<< nsubstratencontact >>
rect -239 72 -235 76
rect -227 72 -223 76
rect -196 72 -192 76
rect -166 72 -162 76
rect -141 72 -137 76
rect -123 72 -119 76
rect -105 72 -101 76
rect -94 72 -90 76
<< labels >>
rlabel metal1 -163 -124 -163 -124 1 Vbias3
rlabel metal1 -237 -11 -237 -11 1 Vbiasp
rlabel metal1 -209 74 -209 74 1 Vdd
rlabel metal1 -200 -188 -200 -188 1 gnd
rlabel metal1 -101 -9 -101 -9 1 Vbias2
rlabel metal1 -118 65 -118 65 1 Vbias1
<< end >>
